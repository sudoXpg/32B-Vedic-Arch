module nop();
    always @(*)
        begin
            #0; 
        end
endmodule
